`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Caldeira & Silva Lda.                                               //
// Engineer: Rui Caldeira, Joel Silva
// 
// Create Date:    15:47:12 04/10/2007 
// Design Name: 
// Module Name:    Multiplication
// Project Name: Calculadora Simples
// Target Devices: 
// Tool versions: 
// Description: M�dulo que multiplica 2 n�meros bin�rios pelo m�todo de Booth.
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Multiplication(mul1,mul2,butMUL,relogio,resMUL);

	input [8:0] mul1; 		//multiplicando
	input [8:0] mul2;			//multiplicador
	input butMUL;				//botao de multiplicacao
	input relogio;
	output [17:0] resMUL;	//resultado de multiplicacao

  	reg [8:0] mu1neg;			//negativo do multiplicando em 2s Complement
	reg [17:0] resMUL;
	reg [18:0] a;				//vector intermedio auxiliar ao calculo pelo metodo de booth
	reg [18:0] s;				//vector intermedio auxiliar ao calculo pelo metodo de booth
	reg [18:0] p;				//vector intermedio auxiliar ao calculo pelo metodo de booth

	reg [18:0] c;				//vectores auxilares 'a soma no metodo de booth
   reg [18:0] d;				//vectores auxilares 'a soma no metodo de booth
	
//variavel intermedia de auxilio ao 2s Complement, 
//toma valor ha1true se ja encontrou o primeiro 1	
	
	parameter ha1true=1'b1;
	parameter ha1false=1'b0;
	
	reg ha1 = ha1false;
	
	parameter state0	= 5'b11111;
	parameter state1  = 5'b00000;
   parameter state2  = 5'b00001;
   parameter state3  = 5'b00010;
   parameter state4  = 5'b00011;
   parameter state5  = 5'b00100;
   parameter state6  = 5'b00101;
   parameter state7  = 5'b00110;
   parameter state8  = 5'b00111;
   parameter state9  = 5'b01000;
	parameter state10 = 5'b01001;
	parameter state11 = 5'b01010;
	parameter state12 = 5'b01011;
	parameter state13 = 5'b01100;
	parameter state14 = 5'b01101;
	parameter state15 = 5'b01110;
	parameter state16 = 5'b01111;
	parameter state17 = 5'b10000;
	parameter state18 = 5'b10001;
	parameter state19 = 5'b10010;
	parameter state20 = 5'b10011;

   reg [3:0] state = state0;	

	always @ (negedge butMUL)		//sempre que o botao multiplicacao e' carregado
	begin

	state = state1;

	end

	always @ (negedge relogio)
	begin

// Nega��o em nota��o Two's Complement --- INICIO ---

        case (state)
            state1 : begin

		mu1neg[0] = mul1[0];
	
		state <=state2;
            end
            state2 : begin
				
		if (mul1[0] == 1'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end
 
		mu1neg[1] = mul1[1] ^ ha1; //xor dos do bit e do ha1

	state <=state3;		
            end
            state3 : begin
				
		if (mul1[1] == 1'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end
 
		mu1neg[2] = mul1[2] ^ ha1; //xor dos do bit e do ha1

	state <=state4;				
            end
            state4 : begin
				
		if (mul1[2] == 1'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end
 
		mu1neg[3] = mul1[3] ^ ha1; //xor dos do bit e do ha1

	state <=state5;		
            end
            state5 : begin
				
		if (mul1[3] == 1'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end
 
		mu1neg[4] = mul1[4] ^ ha1; //xor dos do bit e do ha1

	state <=state6;				
            end
            state6 : begin
				
		if (mul1[4] == 1'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end
 
		mu1neg[5] = mul1[5] ^ ha1; //xor dos do bit e do ha1

	state <=state7;				
            end
            state7 : begin
				
		if (mul1[5] == 1'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end
 
		mu1neg[6] = mul1[6] ^ ha1; //xor dos do bit e do ha1

	state <=state8;				
            end
            state8 : begin
				
		if (mul1[6] == 1'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end
 
		mu1neg[7] = mul1[7] ^ ha1; //xor dos do bit e do ha1

	state <=state9;				
            end
            state9 : begin
				
		if (mul1[7] == 1'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end
 
		mu1neg[8] = mul1[8] ^ ha1; //xor dos do bit e do ha1

	state <=state10;				
        end
		  
				state10 : begin
		
		a = {mul1,9'b000000000,1'b0};
		s = {mu1neg,9'b000000000,1'b0};
		p = {9'b000000000,mul2,1'b0};

	state <=state11;
		  end
		  
				state11 : begin
		
			if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

	state <=state12;
	
			end
			
				state12 : begin
		
			if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

	state <=state13;
	
			end
			
				state13 : begin
		
			if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

	state <=state14;
	
			end

				state14 : begin
		
			if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

	state <=state15;
	
			end

				state15 : begin
		
			if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

	state <=state16;
	
			end
			
				state16 : begin
		
			if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

	state <=state17;
	
			end
			
				state17 : begin
		
			if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

	state <=state18;
	
			end
			
				state18 : begin
		
			if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

	state <=state19;
	
			end

				state19 : begin
		
			if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

	state <=state20;
	
			end
			
			state20 : begin
			
			resMUL = p  >>> 1;
			
			state <=state0;
			end
        
		  endcase

end
endmodule		  
// Nega��o em nota��o Two's Complement --- FIM ---


/*

	always @ (negedge butMUL)		//sempre que o botao e' carregado
	
	begin
	
	ha1 = 0;						
	
// Nega��o em nota��o Two's Complement --- INICIO ---

// O primeiro bit � igual

	mu1neg[0] = mul1[0];

// Verifica se o bit anterior � 1 e se ha1 ainda � 0. Se TRUE, muda valor de ha1 para 1.
	
		if (mul1[0] == 'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end

		mu1neg[1] = mul1[1] ^ ha1;

// Verifica se o bit anterior � 1 e se ha1 ainda � 0. Se TRUE, muda valor de ha1 para 1.
	
		if (mul1[1] == 'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end

		mu1neg[2] = mul1[2] ^ ha1;

// Verifica se o bit anterior � 1 e se ha1 ainda � 0. Se TRUE, muda valor de ha1 para 1.
	
		if (mul1[2] == 'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end

		mu1neg[3] = mul1[3] ^ ha1;

// Verifica se o bit anterior � 1 e se ha1 ainda � 0. Se TRUE, muda valor de ha1 para 1.
	
		if (mul1[3] == 'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end

		mu1neg[4] = mul1[4] ^ ha1;

// Verifica se o bit anterior � 1 e se ha1 ainda � 0. Se TRUE, muda valor de ha1 para 1.
	
		if (mul1[4] == 'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end

		mu1neg[5] = mul1[5] ^ ha1;

// Verifica se o bit anterior � 1 e se ha1 ainda � 0. Se TRUE, muda valor de ha1 para 1.
	
		if (mul1[5] == 'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end

		mu1neg[6] = mul1[6] ^ ha1;

// Verifica se o bit anterior � 1 e se ha1 ainda � 0. Se TRUE, muda valor de ha1 para 1.
	
		if (mul1[6] == 'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end

		mu1neg[7] = mul1[7] ^ ha1;

// Verifica se o bit anterior � 1 e se ha1 ainda � 0. Se TRUE, muda valor de ha1 para 1.
	
		if (mul1[7] == 'b1 & ha1 == ha1false)
		begin
	
		ha1 = ha1true;
		
		end

		mu1neg[8] = mul1[8] ^ ha1;

	
// Nega��o em nota��o Two's Complement --- FIM ---

// Constru��o dos vectores interm�dios para a multiplica��o por Booth

	a = {mul1,9'b000000000,1'b0};
	s = {mu1neg,9'b000000000,1'b0};
	p = {9'b000000000,mul2,1'b0};
	
//	Primeiro passo dos Y passos do Booth (Y = n� de digitos do multiplicador) -- INICIO --
	
	if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

//	Primeiro passso dos Y passos do Booth (Y = n� de digitos do multiplicador) -- FIM --	

if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c  >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c  >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c  >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c  >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c  >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c  >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

if (p[0] ~^ p[1])
   begin
		p = p >>> 1; 
   end
	else
	begin
		if (p[0] == 0 & p[1] == 1)
		begin
			
			
		c[0] = p[0] ^ a[0];
		c[1] = p[1] ^ a[1] ^ p[0] & a[0];
		c[2] = p[2] ^ a[2] ^ a[1] | ~a[1] & p[1] & p[0] & a[0];
		c[3] = p[3] ^ a[3] ^ a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]);
		c[4] = p[4] ^ a[4] ^ a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]));
		c[5] = p[5] ^ a[5] ^ a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])));
		c[6] = p[6] ^ a[6] ^ a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))));
		c[7] = p[7] ^ a[7] ^ a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))));
		c[8] = p[8] ^ a[8] ^ a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))));
		c[9] = p[9] ^ a[9] ^ a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))));
		c[10] = p[10] ^ a[10] ^ a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))));
		c[11] = p[11] ^ a[11] ^ a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))));
		c[12] = p[12] ^ a[12] ^ a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))));
		c[13] = p[13] ^ a[13] ^ a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))));
		c[14] = p[14] ^ a[14] ^ a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))));
		c[15] = p[15] ^ a[15] ^ a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))));
		c[16] = p[16] ^ a[16] ^ a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))));
		c[17] = p[17] ^ a[17] ^ a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0])))))))))))))));
		c[18] = p[18] ^ a[18] ^ a[17] | ~a[17] & p[17] & (a[16] | ~a[16] & p[16] & (a[15] | ~a[15] & p[15] & (a[14] | ~a[14] & p[14] & (a[13] | ~a[13] & p[13] & (a[12] | ~a[12] & p[12] & (a[11] | ~a[11] & p[11] & (a[10] | ~a[10] & p[10] & (a[9] | ~a[9] & p[9] & (a[8] | ~a[8] & p[8] & (a[7] | ~a[7] & p[7] & (a[6] | ~a[6] & p[6] & (a[5] | ~a[5] & p[5] & (a[4] | ~a[4] & p[4] & (a[3] | ~a[3] & p[3] & (a[2] | ~a[2] & p[2] & (a[1] | ~a[1] & p[1] & p[0] & a[0]))))))))))))))));
	
		p = c  >>> 1;
		
		end
		
		else
		begin
		
		d[0] = p[0] ^ s[0];
		d[1] = p[1] ^ s[1] ^ p[0] & s[0];
		d[2] = p[2] ^ s[2] ^ s[1] | ~s[1] & p[1] & p[0] & s[0];
		d[3] = p[3] ^ s[3] ^ s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]);
		d[4] = p[4] ^ s[4] ^ s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]));
		d[5] = p[5] ^ s[5] ^ s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])));
		d[6] = p[6] ^ s[6] ^ s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))));
		d[7] = p[7] ^ s[7] ^ s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))));
		d[8] = p[8] ^ s[8] ^ s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))));
		d[9] = p[9] ^ s[9] ^ s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))));
		d[10] = p[10] ^ s[10] ^ s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))));
		d[11] = p[11] ^ s[11] ^ s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))));
		d[12] = p[12] ^ s[12] ^ s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))));
		d[13] = p[13] ^ s[13] ^ s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))));
		d[14] = p[14] ^ s[14] ^ s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))));
		d[15] = p[15] ^ s[15] ^ s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))));
		d[16] = p[16] ^ s[16] ^ s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))));
		d[17] = p[17] ^ s[17] ^ s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0])))))))))))))));
		d[18] = p[18] ^ s[18] ^ s[17] | ~s[17] & p[17] & (s[16] | ~s[16] & p[16] & (s[15] | ~s[15] & p[15] & (s[14] | ~s[14] & p[14] & (s[13] | ~s[13] & p[13] & (s[12] | ~s[12] & p[12] & (s[11] | ~s[11] & p[11] & (s[10] | ~s[10] & p[10] & (s[9] | ~s[9] & p[9] & (s[8] | ~s[8] & p[8] & (s[7] | ~s[7] & p[7] & (s[6] | ~s[6] & p[6] & (s[5] | ~s[5] & p[5] & (s[4] | ~s[4] & p[4] & (s[3] | ~s[3] & p[3] & (s[2] | ~s[2] & p[2] & (s[1] | ~s[1] & p[1] & p[0] & s[0]))))))))))))))));
	
		p = d  >>> 1;
		
		end
end

//FIM dos Y passos!!!	

// Por fim vamos eliminar o algarismo menos significativo.

     resMUL = p  >>> 1;
	  
end	

*/
	
